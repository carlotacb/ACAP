--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.cte_tipos_deco_camino_pkg.all;

package cte_tipos_deco_camino_ModSecu_pkg is

-- subtipos y constantes utilizadas para el control del camino de datos
-- y operacion en el mismo de una instruccion

constant mSI_relat: st_mSI:= '0';

end package cte_tipos_deco_camino_ModSecu_pkg;

