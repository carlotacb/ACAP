--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_nucleo_pkg is

constant retBRES: time := 14 ns;
constant retBRLE: time := 10 ns;
constant retBRdeco: time := 8 ns;
constant retsuma: time := 16 ns;
constant retreg: time:= 2 ns;
--constant retBCDaDPD: time:= 1 ns;
--constant retDPDaBCD: time:= 1 ns;

end package retardos_nucleo_pkg;

