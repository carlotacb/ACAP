--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_cntl_seg_pkg is

constant retLDRD: time := 1 ns;
constant retLDD: time := 2 ns;
constant retLDRS: time := 1 ns;
constant retLGR: time := 1 ns;

end package retardos_cntl_seg_pkg;

