--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_even_pkg is

constant retexcepMD: time := 1 ns;
constant retexcepMI: time := 1 ns;

constant retlogicaexcep: time := 2 ns;

end package retardos_even_pkg;
