--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_bcd_compresion_pkg is

constant retBCDaDPD: time:= 1 ns;
constant retDPDaBCD: time:= 1 ns;

end package retardos_bcd_compresion_pkg;

