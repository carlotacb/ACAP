--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_cntl_seg_C_pkg is

constant retLDC: time := 1 ns;
constant retLDRD_C: time := 2 ns;

end package retardos_cntl_seg_C_pkg;

