--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_RegDes_pkg is

constant retREGDES: time := 1 ns;

end package retardos_RegDes_pkg;
